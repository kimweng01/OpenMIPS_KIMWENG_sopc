library verilog;
use verilog.vl_types.all;
entity OpenMIPS_KIMWENG_sopc_tb is
end OpenMIPS_KIMWENG_sopc_tb;
