library verilog;
use verilog.vl_types.all;
entity ex is
    port(
        inst_i          : in     vl_logic_vector(31 downto 0);
        aluop_i         : in     vl_logic_vector(7 downto 0);
        alusel_i        : in     vl_logic_vector(2 downto 0);
        reg1_i          : in     vl_logic_vector(31 downto 0);
        reg2_i          : in     vl_logic_vector(31 downto 0);
        wd_i            : in     vl_logic_vector(4 downto 0);
        wreg_i          : in     vl_logic;
        hi_i            : in     vl_logic_vector(31 downto 0);
        lo_i            : in     vl_logic_vector(31 downto 0);
        wb_hi_i         : in     vl_logic_vector(31 downto 0);
        wb_lo_i         : in     vl_logic_vector(31 downto 0);
        wb_whilo_i      : in     vl_logic;
        mem_hi_i        : in     vl_logic_vector(31 downto 0);
        mem_lo_i        : in     vl_logic_vector(31 downto 0);
        mem_whilo_i     : in     vl_logic;
        annul_i         : in     vl_logic;
        maddsub_temp_i  : in     vl_logic_vector(63 downto 0);
        div_temp_i      : in     vl_logic_vector(63 downto 0);
        cnt_mult_i      : in     vl_logic;
        cnt_div_i       : in     vl_logic_vector(4 downto 0);
        link_addr_i     : in     vl_logic_vector(31 downto 0);
        dlyslot_now_i   : in     vl_logic;
        mem_cp0_reg_we  : in     vl_logic;
        mem_cp0_reg_wr_addr: in     vl_logic_vector(4 downto 0);
        mem_cp0_reg_data: in     vl_logic_vector(31 downto 0);
        wb_cp0_reg_we   : in     vl_logic;
        wb_cp0_reg_wr_addr: in     vl_logic_vector(4 downto 0);
        wb_cp0_reg_data : in     vl_logic_vector(31 downto 0);
        cp0_reg_data_i  : in     vl_logic_vector(31 downto 0);
        current_inst_addr_i: in     vl_logic_vector(31 downto 0);
        excepttype_i    : in     vl_logic_vector(31 downto 0);
        wd_o            : out    vl_logic_vector(4 downto 0);
        wreg_o          : out    vl_logic;
        wdata_o         : out    vl_logic_vector(31 downto 0);
        hi_o            : out    vl_logic_vector(31 downto 0);
        lo_o            : out    vl_logic_vector(31 downto 0);
        whilo_o         : out    vl_logic;
        maddsub_temp_o  : out    vl_logic_vector(63 downto 0);
        div_temp_o      : out    vl_logic_vector(63 downto 0);
        cnt_mult_o      : out    vl_logic;
        cnt_div_o       : out    vl_logic_vector(4 downto 0);
        aluop_o         : out    vl_logic_vector(7 downto 0);
        mem_addr_o      : out    vl_logic_vector(31 downto 0);
        reg2_o          : out    vl_logic_vector(31 downto 0);
        cp0_reg_we_o    : out    vl_logic;
        cp0_reg_wr_addr_o: out    vl_logic_vector(4 downto 0);
        cp0_reg_data_o  : out    vl_logic_vector(31 downto 0);
        cp0_reg_rd_addr_o: out    vl_logic_vector(4 downto 0);
        stallreq        : out    vl_logic;
        dlyslot_now_o   : out    vl_logic;
        excepttype_o    : out    vl_logic_vector(31 downto 0);
        current_inst_addr_o: out    vl_logic_vector(31 downto 0)
    );
end ex;
